class test_i2cmb_reg_transactions extends ncsu_component; 
endclass