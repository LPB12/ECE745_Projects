class test_i2cmb_reg_faultaddrs extends ncsu_component; 
endclass