class test_i2cmbFSM_starts extends ncsu_component; 
endclass