class i2c_monitor extends ncsu_component#(.T(i2c_transaction));

  // i2c_configuration configuration;
  // virtual i2c_if bus;

  // T monitored_trans;
  // ncsu_component #(T) agent;

  
endclass
