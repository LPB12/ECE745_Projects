package i2c_pkg;
    import data_pkg::*;
endpackage