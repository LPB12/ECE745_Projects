class test_i2cmbFSM_writefirst extends ncsu_component; 
endclass