class test_i2cmbFSM_stops extends ncsu_component; 
endclass