class wb_coverage extends ncsu_configuration;
  
endclass